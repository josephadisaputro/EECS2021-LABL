module LabL8;

reg signed[31:0] a, b;
reg ctrl;
wire signed[31:0] z;
wire cout;

yArith arith(z, cout, a, b, ctrl);

initial 
begin

		a = 32'b1001;
		b = 32'b1101;
		ctrl = 0;
		#1 $display("a=%b b=%b ctrl=%b z=%b cout=%b", a, b, ctrl, z, cout);
		#1 $display("a=%d b=%d ctrl=%b z=%d cout=%b", a, b, ctrl, z, cout);

end
endmodule
